interface program_counter_interface(input logic CLK_n);
    logic Cp;
    logic Ep;
    logic CLR_n;
    logic [3:0] w_bus_addr;
endinterface