class monitor;
    virtual program_counter_interface pc_if;
    mailbox scb_mbx;


endclass
